; VGA Memory Map 
; .COE file with hex coefficients 
; Height: 16, Width: 16

memory_initialization_radix=2;
memory_initialization_vector=
0001,0001,0001,0001,0001,0001,0001,0001,0001,0001,0001,0001,0001,0001,0001,
0001,0001,0000,0000,0000,0100,0001,1000,0001,0100,0000,0000,0000,0000,0001,
0001,0110,0011,0000,0000,0100,0000,0111,0000,0100,0000,0011,0001,0000,0001,
0001,0001,0000,0000,0011,0100,0000,0000,0000,0100,0011,0110,0011,0000,0001,
0001,0000,0100,0000,0000,0100,0000,0011,0000,0100,0000,0011,0001,0000,0001,
0001,0110,0100,0000,0000,0100,0000,0000,0000,0100,0000,0000,0000,0000,0001,
0001,0000,0100,0000,0000,0100,0000,0000,0000,0100,0000,0000,0000,0000,0001,
0001,0001,0001,0001,0001,0001,0000,0010,0000,0001,0001,0001,0001,0001,0001,
0001,0000,0000,0000,0100,0100,0000,0000,0000,0100,0001,0000,0011,0100,0001,
0001,0000,0011,0100,0100,0100,0000,0000,0000,0100,0001,0000,0100,0110,0001,
0001,0000,0100,0011,0100,0100,0000,0000,0000,0100,0001,0100,0001,0001,0001,
0001,0000,0000,0000,0100,0100,0000,0000,0000,0100,0001,0011,0000,0000,0001,
0001,0000,0100,0000,0100,0100,0000,0000,0110,0100,0000,0000,0001,0000,0001,
0001,0100,0110,0100,0100,0100,0000,0000,0000,0100,0001,0000,0000,0110,0001,
0001,0001,0001,0001,0001,0001,0001,0001,0001,0001,0001,0001,0001,0001,0001,
